library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity flappy_game_top is
    Port (
        CLOCK_50      : in  std_logic;
        RESET_N       : in  std_logic;
        -- PS/2 Mouse
        PS2_CLK       : inout std_logic;
        PS2_DAT       : inout std_logic;
        -- VGA Output
        VGA_R         : out std_logic_vector(3 downto 0);
        VGA_G         : out std_logic_vector(3 downto 0);
        VGA_B         : out std_logic_vector(3 downto 0);
        VGA_HS        : out std_logic;
        VGA_VS        : out std_logic;
        -- Push buttons
        KEY           : in  std_logic_vector(1 downto 0)
    );
end flappy_game_top;

architecture Structural of flappy_game_top is

    signal clk_25mhz     : std_logic;
    signal reset         : std_logic;
    
    -- VGA sync
    signal pixel_row     : std_logic_vector(9 downto 0);
    signal pixel_col     : std_logic_vector(9 downto 0);
    signal video_on      : std_logic;

    -- Mouse output
    signal left_btn      : std_logic;
    signal right_btn     : std_logic;
    signal mouse_x       : std_logic_vector(9 downto 0);
    signal mouse_y       : std_logic_vector(9 downto 0);

    -- Bird display signal
    signal bird_on       : std_logic;
    signal red, green, blue : std_logic;  -- FIXED to single-bit

begin

    reset <= not RESET_N;

    -- Clock divider to 25 MHz
    process(CLOCK_50)
    begin
        if rising_edge(CLOCK_50) then
            clk_25mhz <= not clk_25mhz;
        end if;
    end process;

    -- VGA controller
    vga_sync_inst : entity work.VGA_SYNC
        port map (
            clock_25Mhz      => clk_25mhz,
            red              => red,
            green            => green,
            blue             => blue,
            red_out          => VGA_R(0),
            green_out        => VGA_G(0),
            blue_out         => VGA_B(0),
            horiz_sync_out   => VGA_HS,
            vert_sync_out    => VGA_VS,
            pixel_row        => pixel_row,
            pixel_column     => pixel_col
        );

    -- PS/2 mouse interface
    mouse_inst : entity work.MOUSE
        port map (
            clock_25Mhz         => clk_25mhz,
            reset               => reset,
            mouse_data          => PS2_DAT,
            mouse_clk           => PS2_CLK,
            left_button         => left_btn,
            right_button        => right_btn,
            mouse_cursor_row    => mouse_y,
            mouse_cursor_column => mouse_x
        );

    -- Bird logic: treat the bird like a bouncing ball for now
    ball_inst : entity work.bouncy_ball
        port map (
            clk        => clk_25mhz,
            reset      => reset,
            click      => left_btn,
            pixel_row  => pixel_row,
            pixel_col  => pixel_col,
            bird_on    => bird_on
        );

    -- Yellow bird: Red + Green on, Blue off
    red   <= bird_on;
    green <= bird_on;
    blue  <= '0';

    -- Replicate single-bit color over 4-bit VGA outputs
    VGA_R <= (others => red)   when video_on = '1' else (others => '0');
    VGA_G <= (others => green) when video_on = '1' else (others => '0');
    VGA_B <= (others => blue)  when video_on = '1' else (others => '0');

end Structural;

