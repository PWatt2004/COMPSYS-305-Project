LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
ENTITY flappy_bird_base IS
    PORT (
        CLOCK_50 : IN STD_LOGIC; -- 50 MHz input clock signal, drives the entire system for timing and synchronization.
        RESET_N : IN STD_LOGIC; -- Active-low reset signal; logic '0' resets the system to initial state.
        PS2_CLK : INOUT STD_LOGIC; -- PS/2 keyboard clock line (bidirectional). The PS2_CLK signal synchronizes data transmission for PS/2 devices (keyboard), ensuring each data bit from PS2_DAT is sampled correctly on clock edges. Often, devices hold the clock low to signal start of communication.
        PS2_DAT : INOUT STD_LOGIC; -- PS/2 keyboard data line (bidirectional). Carries serial data between the keyboard and FPGA. Bits are sent synchronously with PS2_CLK, including start, data, parity, and stop bits, allowing key press/release codes to be received and processed by the game.
        VGA_R : OUT STD_LOGIC_VECTOR(3 DOWNTO 0); -- Red color channel output (4-bit) for VGA display. For each pixel clock cycle, these 4 bits determine the red intensity (0-15 levels). Together with VGA_G and VGA_B, this defines the pixel's final RGB color. The current pixel location is determined by sync signals and internal counters.
        VGA_G : OUT STD_LOGIC_VECTOR(3 DOWNTO 0); -- Green color channel output (4-bit) for VGA display. Similar to VGA_R, it defines green intensity per pixel (0-15 levels). The combination of VGA_R, VGA_G, VGA_B for each pixel clock updates the screen's color at that pixel coordinate.
        VGA_B : OUT STD_LOGIC_VECTOR(3 DOWNTO 0); -- Blue color channel output (4-bit) for VGA display. Controls blue intensity (0-15 levels) per pixel. During active video time, the FPGA updates VGA_B (along with R and G) on each pixel clock to paint the screen with desired colors (bird, pipes, background).
        VGA_HS : OUT STD_LOGIC; -- Horizontal sync pulse for VGA. Generated by the FPGA at specific intervals to signal the end of a horizontal scanline. When VGA_HS pulses low, the display circuitry knows to reset the horizontal pixel counter and move to the next line. It helps align the timing of pixel data (R,G,B) to the screen's scanline refresh.
        VGA_VS : OUT STD_LOGIC; -- Vertical sync pulse for VGA. Pulses low once per screen frame to signal the end of vertical scanning. It resets the vertical pixel counter and starts a new frame refresh. VGA_VS combined with VGA_HS ensures the monitor knows when to start drawing from (0,0) again, maintaining correct image placement and timing.
        LEDR : OUT STD_LOGIC_VECTOR(9 DOWNTO 0); -- 10-bit output for LEDs; each bit controls one LED (1=on, 0=off).
        SW : IN STD_LOGIC_VECTOR(9 DOWNTO 0); -- 10-bit input from switches; each bit reflects a switch state (1=on, 0=off).
        HEX0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0); -- 7-segment output for HEX0 display; controls segments a-g (1=on, 0=off).
        HEX1 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0); -- 7-segment output for HEX1 display; controls segments a-g (1=on, 0=off).
        HEX2 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0) -- 7-segment output for HEX2 display; controls segments a-g (1=on, 0=off).
    );
END flappy_bird_base;
ARCHITECTURE top OF flappy_bird_base IS --Defines the behavior of this top-level component

    -- The char_rom component is used to retrieve font data for rendering characters on the screen.
    -- It acts as a read-only memory (ROM) that stores the pixel patterns for each character in a font set.
    -- Each character is represented as a 5x7 pixel grid, and the ROM outputs the corresponding pixel value.

    COMPONENT char_rom
        PORT (
            character_address : IN STD_LOGIC_VECTOR(5 DOWNTO 0); -- Input address specifying which character's font data to retrieve (6 bits, allowing for 64 characters).
            font_row : IN STD_LOGIC_VECTOR(2 DOWNTO 0); -- Input specifying the row of the character's pixel grid (3 bits, allowing for 8 rows).
            font_col : IN STD_LOGIC_VECTOR(2 DOWNTO 0); -- Input specifying the column of the character's pixel grid (3 bits, allowing for 8 columns).
            clock : IN STD_LOGIC; -- Clock signal to synchronize the ROM read operation.
            rom_mux_output : OUT STD_LOGIC -- Output signal providing the pixel value (1=on, 0=off) for the specified character, row, and column.
        );
    END COMPONENT;

    -- Declare a component named "background" that will be instantiated in the architecture.
    COMPONENT background
        PORT (
            clk : IN STD_LOGIC; -- Input clock signal to synchronize the background rendering logic.
            pixel_row : IN STD_LOGIC_VECTOR(9 DOWNTO 0); -- Input specifying the current pixel row (10-bit vector, supports up to 1024 rows).
            pixel_column : IN STD_LOGIC_VECTOR(9 DOWNTO 0); -- Input specifying the current pixel column (10-bit vector, supports up to 1024 columns).
            bg_red : OUT STD_LOGIC; -- Output signal for the red color channel of the background (1-bit, on/off).
            bg_green : OUT STD_LOGIC; -- Output signal for the green color channel of the background (1-bit, on/off).
            bg_blue : OUT STD_LOGIC -- Output signal for the blue color channel of the background (1-bit, on/off).
        );
    END COMPONENT;

    -- Declare a component named "display_text" that will be instantiated in the architecture.
    COMPONENT display_text
        PORT (
            clk : IN STD_LOGIC; -- Input clock signal to synchronize the text rendering logic.
            pixel_row : IN STD_LOGIC_VECTOR(9 DOWNTO 0); -- Input specifying the current pixel row (10-bit vector, supports up to 1024 rows).
            pixel_column : IN STD_LOGIC_VECTOR(9 DOWNTO 0); -- Input specifying the current pixel column (10-bit vector, supports up to 1024 columns).
            score : IN STD_LOGIC_VECTOR(11 DOWNTO 0); -- Input signal representing the player's score (12-bit vector, supports values up to 4095).
            health_percentage : IN STD_LOGIC_VECTOR(11 DOWNTO 0); -- Input signal representing the player's health percentage (12-bit vector, supports values up to 4095).
            text_rgb : OUT STD_LOGIC_VECTOR(11 DOWNTO 0); -- Output signal for the RGB color of the text (12-bit vector, 4 bits per color channel).
            text_on : OUT STD_LOGIC -- Output signal indicating whether the text is currently being displayed (1 = on, 0 = off).
        );
    END COMPONENT;

    -- Type definition: an unconstrained array of integers, used for collections like pipe positions.
    TYPE INTEGER_VECTOR IS ARRAY (NATURAL RANGE <>) OF INTEGER;
    -- 25 MHz clock signal for VGA timing. Derived from main 50 MHz clock by dividing by 2. Drives pixel scanning.
    SIGNAL clk_25 : STD_LOGIC;
    -- Single-bit outputs controlling the current pixel's red, green, and blue states on VGA. These are updated each pixel clock.
    SIGNAL red, green, blue : STD_LOGIC;
    -- Current pixel's vertical (row) and horizontal (column) position on the screen (0 to 639 columns, 0 to 479 rows). Used to determine what should be drawn at each pixel.
    SIGNAL pixel_row, pixel_column : STD_LOGIC_VECTOR(9 DOWNTO 0);
    -- Mouse cursor position on screen. Updated from PS/2 mouse input. Used for interactive controls (menus, maybe aiming or flapping).
    SIGNAL mouse_row, mouse_col : STD_LOGIC_VECTOR(9 DOWNTO 0);
    -- Mouse button states. '1' if pressed. Can be used for bird flapping (left_button) or other actions (right_button).
    SIGNAL left_button, right_button : STD_LOGIC;
    -- Bird's vertical position in pixels. Controls where the bird is drawn on screen (Y coordinate).
    SIGNAL bird_y : INTEGER;
    -- Bird's current vertical velocity. Positive values move the bird down, negative values up. Updated by gravity and flap inputs.
    SIGNAL bird_velocity : INTEGER;
    -- Collision detection signal. '1' when bird collides with a pipe. Triggers game over or health reduction.
    SIGNAL pipe_hit : STD_LOGIC;
    -- Array holding X positions of up to 4 pipes. Controls where pipes are drawn horizontally on screen.
    SIGNAL pipe_x_array : INTEGER_VECTOR(0 TO 3);
    -- Flattened output of pipe X positions for driving VGA output logic. Combines multiple pipes into a single bus.
    SIGNAL pipe_x_out : STD_LOGIC_VECTOR(39 DOWNTO 0);
    -- Flattened output of pipe Y positions (vertical gaps). Controls pipe hole placement for VGA drawing.
    SIGNAL pipe_y_out : STD_LOGIC_VECTOR(39 DOWNTO 0);
    -- Array holding Y positions of up to 4 pipes (typically the top edge of the gap). Used for collision and rendering.
    SIGNAL pipe_y_array : INTEGER_VECTOR(0 TO 3);
    -- Internal signal mirroring VGA vertical sync. Used for frame updates and synchronizing game logic with display refresh.
    SIGNAL vsync_internal : STD_LOGIC;
    -- Background color signals for red, green, and blue channels. Determines what background color is shown at each pixel location.
    SIGNAL bg_red, bg_green, bg_blue : STD_LOGIC;
    -- Current score represented in BCD or raw binary (12-bit wide). Drives score display on 7-segment or on-screen text.
    SIGNAL score : STD_LOGIC_VECTOR(11 DOWNTO 0) := (OTHERS => '0');
    -- Bird's health represented as a percentage (0-100%) in a 12-bit vector. Drives health bar or UI display.
    SIGNAL health_percentage : STD_LOGIC_VECTOR(11 DOWNTO 0) := (OTHERS => '1');
    -- RGB signal used for displaying text on screen. 12-bit (likely 4-bit per color channel). Drives pixel color when text is rendered.
    SIGNAL text_rgb_signal : STD_LOGIC_VECTOR(11 DOWNTO 0);
    -- Text rendering flag. '1' when current pixel overlaps with a text glyph (e.g., score numbers). Used to decide whether to draw text or game graphics.
    SIGNAL text_on_signal : STD_LOGIC;
    -- Constant horizontal position for the bird (X coordinate). The bird stays at this X position; only Y changes to simulate movement.
    CONSTANT bird_x : INTEGER := 100;
    -- Used for dividing or positioning, often related to screen boundaries or object placement. Here, 590 might represent bottom ground level (screen height - ground height).
    SIGNAL number : INTEGER := 590;
    -- Binary-coded decimal outputs for hundreds, tens, and ones digits. Drives 7-segment displays or on-screen numeric rendering.
    SIGNAL hundreds, tens, ones : STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN
    -- Instantiate 7-segment decoders
    hundred_display : ENTITY work.BCD_to_SevenSeg
        PORT MAP(
            BCD_digit => hundreds,
            SevenSeg_out => HEX2
        );

    ten_display : ENTITY work.BCD_to_SevenSeg
        PORT MAP(
            BCD_digit => tens,
            SevenSeg_out => HEX1
        );

    one_display : ENTITY work.BCD_to_SevenSeg
        PORT MAP(
            BCD_digit => ones,
            SevenSeg_out => HEX0
        );
    digit_split : PROCESS (number)
        VARIABLE temp : INTEGER;
    BEGIN
        temp := number;
        hundreds <= STD_LOGIC_VECTOR(to_unsigned((temp / 100) MOD 10, 4));
        tens <= STD_LOGIC_VECTOR(to_unsigned((temp / 10) MOD 10, 4));
        ones <= STD_LOGIC_VECTOR(to_unsigned(temp MOD 10, 4));
    END PROCESS digit_split;

    LEDR(0) <= left_button;

    VGA_VS <= vsync_internal;

    clk_divider : PROCESS (CLOCK_50)
        VARIABLE counter : STD_LOGIC := '0';
    BEGIN
        IF rising_edge(CLOCK_50) THEN
            counter := NOT counter;
            clk_25 <= counter;
        END IF;
    END PROCESS;

    vga_inst : ENTITY work.vga_sync
        PORT MAP(
            -- 25 MHz pixel clock input for VGA timing. Drives the pixel scanning logic inside vga_sync.
            -- This ensures that pixels are updated at the correct rate for a 640x480 @ 60Hz VGA display.
            clock_25Mhz => clk_25,
            -- Single-bit red color signal from game logic (e.g., bird, pipes, background).
            -- This is the "raw" red signal deciding whether this current pixel should be red (1) or not (0).
            red => red,
            -- Single-bit green color signal from game logic.
            -- Similar to red, this controls whether the current pixel should have green component active.
            green => green,
            -- Single-bit blue color signal from game logic.
            -- Determines if the blue component is active for the current pixel.
            blue => blue,
            -- Output: drives the 4th bit (MSB) of the VGA red channel.
            -- This maps the internal red signal to the visible VGA output.
            -- Since VGA_R is a 4-bit vector, only bit 3 is used here for simplicity (on/off style graphics).
            red_out => VGA_R(3),
            -- Output: drives the 4th bit (MSB) of the VGA green channel.
            -- Same idea as red_out, this updates VGA_G(3) according to internal green signal.
            green_out => VGA_G(3),
            -- Output: drives the 4th bit (MSB) of the VGA blue channel.
            -- Controls VGA_B(3) based on the internal blue signal, affecting pixel color intensity.
            blue_out => VGA_B(3),
            -- Output: horizontal sync pulse for VGA.
            -- Pulses low at the end of each scanline to signal horizontal retrace.
            -- Tells the monitor to reset its horizontal drawing position.
            horiz_sync_out => VGA_HS,
            -- Output: vertical sync pulse for VGA.
            -- Goes low at the end of a full screen refresh (all lines drawn).
            -- Synchronizes frame redraws and triggers end-of-frame logic.
            -- This is wired to an internal vsync signal for additional game logic use.
            vert_sync_out => vsync_internal,
            -- Output: current pixel row number (Y coordinate, 0-479).
            -- Increments with every completed scanline.
            -- Used by game logic to decide if objects like bird, pipes, background should be drawn at this row.
            pixel_row => pixel_row,
            -- Output: current pixel column number (X coordinate, 0-639).
            -- Increments every pixel clock tick across the screen width.
            -- Helps in deciding horizontal placement of objects (pipes, text, bird sprite, etc.).
            pixel_column => pixel_column
        );
    mouse_inst : ENTITY work.mouse
        PORT MAP(
            clock_25Mhz => clk_25,
            reset => NOT RESET_N,
            mouse_data => PS2_DAT,
            mouse_clk => PS2_CLK,
            left_button => left_button,
            right_button => right_button,
            mouse_cursor_row => mouse_row,
            mouse_cursor_column => mouse_col
        );

    bird_inst : ENTITY work.bird_controller
        PORT MAP(
            clk => vsync_internal,
            reset => NOT RESET_N,
            flap_button => left_button,
            bird_y => bird_y,
            bird_velocity => bird_velocity,
            bird_altitude => number
        );

    background_inst : ENTITY work.background
        PORT MAP(
            clk => clk_25,
            pixel_row => pixel_row,
            pixel_column => pixel_column,
            bg_red => bg_red,
            bg_green => bg_green,
            bg_blue => bg_blue
        );

    pipe_ctrl_inst : ENTITY work.pipe_controller
        PORT MAP(
            clk => vsync_internal,
            reset => NOT RESET_N,
            bird_x => bird_x,
            bird_y => bird_y,
            pipe_hit => pipe_hit,
            pipe_x_out => pipe_x_out,
            pipe_y_out => pipe_y_out
        );

    display_text_inst : ENTITY work.display_text
        PORT MAP(
            clk => clk_25,
            pixel_row => pixel_row,
            pixel_column => pixel_column,
            score => score,
            health_percentage => health_percentage,
            text_rgb => text_rgb_signal,
            text_on => text_on_signal,
            title_on => SW(0),
            score_on => SW(1),
            hp_on => SW(2)
        );

    -- Extract the X positions of pipes from the packed 40-bit pipe_x_out bus.
    -- Each pipe's X coordinate is stored in 10 bits (0-639 range for screen width).
    pipe_x_array(0) <= to_integer(unsigned(pipe_x_out(9 DOWNTO 0))); -- Pipe 0's horizontal position.
    pipe_x_array(1) <= to_integer(unsigned(pipe_x_out(19 DOWNTO 10))); -- Pipe 1's horizontal position.
    pipe_x_array(2) <= to_integer(unsigned(pipe_x_out(29 DOWNTO 20))); -- Pipe 2's horizontal position.
    pipe_x_array(3) <= to_integer(unsigned(pipe_x_out(39 DOWNTO 30))); -- Pipe 3's horizontal position.
    -- Extract the Y positions of pipes (gap top edge) from the packed 40-bit pipe_y_out bus.
    -- Same structure: each pipe's Y coordinate is stored in 10 bits (0-479 range for screen height).
    pipe_y_array(0) <= to_integer(unsigned(pipe_y_out(9 DOWNTO 0))); -- Pipe 0's vertical gap position.
    pipe_y_array(1) <= to_integer(unsigned(pipe_y_out(19 DOWNTO 10))); -- Pipe 1's vertical gap position.
    pipe_y_array(2) <= to_integer(unsigned(pipe_y_out(29 DOWNTO 20))); -- Pipe 2's vertical gap position.
    pipe_y_array(3) <= to_integer(unsigned(pipe_y_out(39 DOWNTO 30))); -- Pipe 3's vertical gap position.
    draw_logic : PROCESS (pixel_row, pixel_column)
        VARIABLE size : INTEGER := 6; -- Defines half-size of bird hitbox for rendering (bird is 12x12 pixels).
    BEGIN

        -- Start by setting the pixel color to the background color by default.
        red <= bg_red;
        green <= bg_green;
        blue <= bg_blue;
        FOR i IN 0 TO 3 LOOP --draw pipes
            IF (to_integer(unsigned(pixel_column)) >= pipe_x_array(i) AND
                to_integer(unsigned(pixel_column)) < pipe_x_array(i) + 20 AND
                (to_integer(unsigned(pixel_row)) < pipe_y_array(i) OR
                to_integer(unsigned(pixel_row)) > pipe_y_array(i) + 100)) THEN

            END IF;
        END LOOP;

        IF ABS(to_integer(unsigned(pixel_column)) - bird_x) < size AND -- draw vird
            ABS(to_integer(unsigned(pixel_row)) - bird_y) < size THEN

            red <= '1';
            green <= '1';
            blue <= '0';
        END IF;

        IF text_on_signal = '1' THEN --draw text
            red <= text_rgb_signal(11); -- Extract red component from text RGB signal.
            green <= text_rgb_signal(5); -- Extract green component.
            blue <= text_rgb_signal(0); -- Extract blue component.
        END IF;

    END PROCESS;

    VGA_R(2 DOWNTO 0) <= (OTHERS => '0'); -- Zero out lower 3 bits of VGA red output.
    VGA_G(2 DOWNTO 0) <= (OTHERS => '0'); -- Zero out lower 3 bits of VGA green output.
    VGA_B(2 DOWNTO 0) <= (OTHERS => '0'); -- Zero out lower 3 bits of VGA blue output.
END top;